//SEQR file
//
class pcie_seqr extends uvm_sequencer#(pcie_tx);
	`uvm_component_utils(pcie_seqr)
	`NEW_COMP
endclass
