import uvm_pkg::*;

module tb_top;
	





	initial begin

		//`uvm_info("TB_TOP","THIS IS IN TOP OF TB",UVM_INFO)
		$display("THSI\n");
	end


endmodule
