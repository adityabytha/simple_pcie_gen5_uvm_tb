//PACKAGE FILE
//includes all files in testbench as a consolidated package
//

package pcie_pkg;
	`include "uvm_commons.sv"
	`include "pcie_env.sv"
	`include "pcie_test_lib.sv"

endpackage
