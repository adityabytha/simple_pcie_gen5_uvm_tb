//PACKAGE FILE
//includes all files in testbench as a consolidated package
//

package pcie_pkg;
	`include "uvm_pkg.sv"
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	//`include "pcie_tl_src.sv"
	//`include "uvm_commons.sv"
	//`include "pcie_env.sv"
	//`include "pcie_test_lib.sv"
	//`include "pcie_tx.sv"



endpackage
