//SEQR file
//
class pcie_seqr extends uvm_sequencer#(uvm_sequence_item);
	`uvm_component_utils(pcie_seqr)
	`NEW_COMP
endclass
/*
class pcie_cpl_seqr extends uvm_sequencer#(pcie_cpl_tx);
	`uvm_component_utils(pcie_cpl_seqr)
	`NEW_COMP
endclass
*/
